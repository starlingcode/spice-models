* C:\Arquivos de Programas\LTC\SwCADIII\lib\sub\regulators.lib


* LM7805 model. 
* No need to use .inc - I've set the .asy symbol to remove the need for .inc.
* (I used the symbol of LT1084, just replaced the LT1084 by LMxxxx and LTC.LIB by regulators.lib) 

.SUBCKT LM7805  1    2    3
* In GND Out
QT6          23  10  2   Q_NPN 0.1
QT7          5   4   10  Q_NPN 0.1
QT5          7   6   5   Q_NPN 0.1
QT1          1   9   8   Q_NPN 0.1
QT3          11  8   7   Q_NPN 0.1
QT2          11  13  12  Q_NPN 0.1
QT17         1   15  14  Q_NPN 10
C2           10  23      4P
R16          12  5       500
R12          16  2       12.1K
QT18         17  23  16  Q_NPN 0.1
D1           18  19  	 D_D 
R11          20  21      850
R5           22  3       100
QT14         24  18  2   Q_NPN 0.1
R21          6   2       2.67K
R20          3   6       640
DZ2          25  26      D_5V1 
R19          1   26      16K
R18          14  3       250M
R17          25  14      380
R15          25  15      1.62K
QT16         1   20  15  Q_NPN 1
QT15         2   24  21  Q_PNP 0.1
*OFF
R14          21  24      4K
C1           27  24      20P
R13          19  2       4K
QT13         24  27  18  Q_NPN 0.1
QT12         20  25  22  Q_NPN 1 
*OFF
QT11         20  28  2   Q_NPN 0.1
*OFF
QT10         20  11  1   Q_PNP 0.1
R10          17  27      16.5K
R9           5   4       1.9K
R8           4   23      26
R7           10  2       1.2K
R6           29  2       1K
QT9          11  11  1   Q_PNP 0.1
QT8          27  16  29  Q_NPN 0.1
QT4          15  6   17  Q_NPN 0.1
DZ1          2   9       D_5V6
R4           1   9       80K
R3           28  2       830
R2           13  28      4.97K
R1           8   13      7K

.MODEL D_5V1 D( IS=10F N=1.16 BV=5.1 IBV=0.5M CJ0 = 1P TT = 10p )
.MODEL D_5V6 D( IS=10F N=1.16 BV=5.6 IBV=5U CJ0 = 1P TT = 10p )
.MODEL Q_NPN NPN( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+       TF=10P TR=1N )
.MODEL Q_PNP PNP( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+      TF=10P TR=1N )
.MODEL D_D D( IS=1F N=1.16 CJ0 = 1P TT = 10p )

.ENDS LM7805

* Pinouts are the same as 7805.

.SUBCKT LM7806  1    2    3
QT6          23  10  2   Q_NPN 0.1
QT7          5   4   10  Q_NPN 0.1
QT5          7   6   5   Q_NPN 0.1
QT1          1   9   8   Q_NPN 0.1
QT3          11  8   7   Q_NPN 0.1
QT2          11  13  12  Q_NPN 0.1
QT17         1   15  14  Q_NPN 10
C2           10  23      4P
R16          12  5       500
R12          16  2       12.1K
QT18         17  23  16  Q_NPN 0.1
D1           18  19  	 D_D 
R11          20  21      850
R5           22  3       100
QT14         24  18  2   Q_NPN 0.1
R21          6   2       2.67K
R20          3   6       1.294K
DZ2          25  26      D_5V1 
R19          1   26      16K
R18          14  3       250M
R17          25  14      380
R15          25  15      1.62K
QT16         1   20  15  Q_NPN 1
QT15         2   24  21  Q_PNP 0.1 
*OFF
R14          21  24      4K
C1           27  24      20P
R13          19  2       4K
QT13         24  27  18  Q_NPN 0.1
QT12         20  25  22  Q_NPN 1 
*OFF
QT11         20  28  2   Q_NPN 0.1
*OFF
QT10         20  11  1   Q_PNP 0.1
R10          17  27      16.5K
R9           5   4       1.9K
R8           4   23      26
R7           10  2       1.2K
R6           29  2       1K
QT9          11  11  1   Q_PNP 0.1
QT8          27  16  29  Q_NPN 0.1
QT4          15  6   17  Q_NPN 0.1
DZ1          2   9       D_5V6
R4           1   9       80K
R3           28  2       830
R2           13  28      4.97K
R1           8   13      7K

.MODEL D_5V1 D( IS=10F N=1.16 BV=5.1 IBV=0.5M CJ0 = 1P TT = 10p )
.MODEL D_5V6 D( IS=10F N=1.16 BV=5.6 IBV=5U CJ0 = 1P TT = 10p )
.MODEL Q_NPN NPN( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+       TF=10P TR=1N )
.MODEL Q_PNP PNP( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+      TF=10P TR=1N )
.MODEL D_D D( IS=1F N=1.16 CJ0 = 1P TT = 10p )

.ENDS LM7806

* Pinouts are the same as 7805.

* Pinouts are the same as 7805.

.SUBCKT LM7808  1    2    3
QT6          23  10  2   Q_NPN 0.1
QT7          5   4   10  Q_NPN 0.1
QT5          7   6   5   Q_NPN 0.1
QT1          1   9   8   Q_NPN 0.1
QT3          11  8   7   Q_NPN 0.1
QT2          11  13  12  Q_NPN 0.1
QT17         1   15  14  Q_NPN 10
C2           10  23      4P
R16          12  5       500
R12          16  2       12.1K
QT18         17  23  16  Q_NPN 0.1
D1           18  19  	 D_D 
R11          20  21      850
R5           22  3       100
QT14         24  18  2   Q_NPN 0.1
R21          6   2       2.67K
R20          3   6       2.60K
DZ2          25  26      D_5V1 
R19          1   26      16K
R18          14  3       250M
R17          25  14      380
R15          25  15      1.62K
QT16         1   20  15  Q_NPN 1
QT15         2   24  21  Q_PNP 0.1 
*OFF
R14          21  24      4K
C1           27  24      20P
R13          19  2       4K
QT13         24  27  18  Q_NPN 0.1
QT12         20  25  22  Q_NPN 1 
*OFF
QT11         20  28  2   Q_NPN 0.1
*OFF
QT10         20  11  1   Q_PNP 0.1
R10          17  27      16.5K
R9           5   4       1.9K
R8           4   23      26
R7           10  2       1.2K
R6           29  2       1K
QT9          11  11  1   Q_PNP 0.1
QT8          27  16  29  Q_NPN 0.1
QT4          15  6   17  Q_NPN 0.1
DZ1          2   9       D_5V6
R4           1   9       80K
R3           28  2       830
R2           13  28      4.97K
R1           8   13      7K

.MODEL D_5V1 D( IS=10F N=1.16 BV=5.1 IBV=0.5M CJ0 = 1P TT = 10p )
.MODEL D_5V6 D( IS=10F N=1.16 BV=5.6 IBV=5U CJ0 = 1P TT = 10p )
.MODEL Q_NPN NPN( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+       TF=10P TR=1N )
.MODEL Q_PNP PNP( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+      TF=10P TR=1N )
.MODEL D_D D( IS=1F N=1.16 CJ0 = 1P TT = 10p )

.ENDS LM7808

.SUBCKT LM7809  1    2    3
QT6          23  10  2   Q_NPN 0.1
QT7          5   4   10  Q_NPN 0.1
QT5          7   6   5   Q_NPN 0.1
QT1          1   9   8   Q_NPN 0.1
QT3          11  8   7   Q_NPN 0.1
QT2          11  13  12  Q_NPN 0.1
QT17         1   15  14  Q_NPN 10
C2           10  23      4P
R16          12  5       500
R12          16  2       12.1K
QT18         17  23  16  Q_NPN 0.1
D1           18  19  	 D_D 
R11          20  21      850
R5           22  3       100
QT14         24  18  2   Q_NPN 0.1
R21          6   2       2.67K
R20          3   6       3.256K
DZ2          25  26      D_5V1 
R19          1   26      16K
R18          14  3       250M
R17          25  14      380
R15          25  15      1.62K
QT16         1   20  15  Q_NPN 1
QT15         2   24  21  Q_PNP 0.1 
*OFF
R14          21  24      4K
C1           27  24      20P
R13          19  2       4K
QT13         24  27  18  Q_NPN 0.1
QT12         20  25  22  Q_NPN 1 
*OFF
QT11         20  28  2   Q_NPN 0.1
*OFF
QT10         20  11  1   Q_PNP 0.1
R10          17  27      16.5K
R9           5   4       1.9K
R8           4   23      26
R7           10  2       1.2K
R6           29  2       1K
QT9          11  11  1   Q_PNP 0.1
QT8          27  16  29  Q_NPN 0.1
QT4          15  6   17  Q_NPN 0.1
DZ1          2   9       D_5V6
R4           1   9       80K
R3           28  2       830
R2           13  28      4.97K
R1           8   13      7K

.MODEL D_5V1 D( IS=10F N=1.16 BV=5.1 IBV=0.5M CJ0 = 1P TT = 10p )
.MODEL D_5V6 D( IS=10F N=1.16 BV=5.6 IBV=5U CJ0 = 1P TT = 10p )
.MODEL Q_NPN NPN( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+       TF=10P TR=1N )
.MODEL Q_PNP PNP( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+      TF=10P TR=1N )
.MODEL D_D D( IS=1F N=1.16 CJ0 = 1P TT = 10p )

.ENDS LM7809

* Pinouts are the same as 7805.

.SUBCKT LM7812  1    2    3
QT6          23  10  2   Q_NPN 0.1
QT7          5   4   10  Q_NPN 0.1
QT5          7   6   5   Q_NPN 0.1
QT1          1   9   8   Q_NPN 0.1
QT3          11  8   7   Q_NPN 0.1
QT2          11  13  12  Q_NPN 0.1
QT17         1   15  14  Q_NPN 10
C2           10  23      4P
R16          12  5       500
R12          16  2       12.1K
QT18         17  23  16  Q_NPN 0.1
D1           18  19  	 D_D 
R11          20  21      850
R5           22  3       100
QT14         24  18  2   Q_NPN 0.1
R21          6   2       2.67K
R20          3   6       5.22K
DZ2          25  26      D_5V1 
R19          1   26      16K
R18          14  3       250M
R17          25  14      380
R15          25  15      1.62K
QT16         1   20  15  Q_NPN 1
QT15         2   24  21  Q_PNP 0.1 
*OFF
R14          21  24      4K
C1           27  24      20P
R13          19  2       4K
QT13         24  27  18  Q_NPN 0.1
QT12         20  25  22  Q_NPN 1 
*OFF
QT11         20  28  2   Q_NPN 0.1
*OFF
QT10         20  11  1   Q_PNP 0.1
R10          17  27      16.5K
R9           5   4       1.9K
R8           4   23      26
R7           10  2       1.2K
R6           29  2       1K
QT9          11  11  1   Q_PNP 0.1
QT8          27  16  29  Q_NPN 0.1
QT4          15  6   17  Q_NPN 0.1
DZ1          2   9       D_5V6
R4           1   9       80K
R3           28  2       830
R2           13  28      4.97K
R1           8   13      7K

.MODEL D_5V1 D( IS=10F N=1.16 BV=5.1 IBV=0.5M CJ0 = 1P TT = 10p )
.MODEL D_5V6 D( IS=10F N=1.16 BV=5.6 IBV=5U CJ0 = 1P TT = 10p )
.MODEL Q_NPN NPN( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+       TF=10P TR=1N )
.MODEL Q_PNP PNP( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+      TF=10P TR=1N )
.MODEL D_D D( IS=1F N=1.16 CJ0 = 1P TT = 10p )

.ENDS LM7812

* Pinouts are the same as '05

.SUBCKT LM7815  1    2    3
QT6          23  10  2   Q_NPN 0.1
QT7          5   4   10  Q_NPN 0.1
QT5          7   6   5   Q_NPN 0.1
QT1          1   9   8   Q_NPN 0.1
QT3          11  8   7   Q_NPN 0.1
QT2          11  13  12  Q_NPN 0.1
QT17         1   15  14  Q_NPN 10
C2           10  23      4P
R16          12  5       500
R12          16  2       12.1K
QT18         17  23  16  Q_NPN 0.1
D1           18  19  	 D_D 
R11          20  21      850
R5           22  3       100
QT14         24  18  2   Q_NPN 0.1
R21          6   2       2.67K
R20          3   6       7.18K
DZ2          25  26      D_5V1 
R19          1   26      16K
R18          14  3       250M
R17          25  14      380
R15          25  15      1.62K
QT16         1   20  15  Q_NPN 1
QT15         2   24  21  Q_PNP 0.1 
*OFF
R14          21  24      4K
C1           27  24      20P
R13          19  2       4K
QT13         24  27  18  Q_NPN 0.1
QT12         20  25  22  Q_NPN 1 
*OFF
QT11         20  28  2   Q_NPN 0.1
*OFF
QT10         20  11  1   Q_PNP 0.1
R10          17  27      16.5K
R9           5   4       1.9K
R8           4   23      26
R7           10  2       1.2K
R6           29  2       1K
QT9          11  11  1   Q_PNP 0.1
QT8          27  16  29  Q_NPN 0.1
QT4          15  6   17  Q_NPN 0.1
DZ1          2   9       D_5V6
R4           1   9       80K
R3           28  2       830
R2           13  28      4.97K
R1           8   13      7K

.MODEL D_5V1 D( IS=10F N=1.16 BV=5.1 IBV=0.5M CJ0 = 1P TT = 10p )
.MODEL D_5V6 D( IS=10F N=1.16 BV=5.6 IBV=5U CJ0 = 1P TT = 10p )
.MODEL Q_NPN NPN( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+       TF=10P TR=1N )
.MODEL Q_PNP PNP( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+      TF=10P TR=1N )
.MODEL D_D D( IS=1F N=1.16 CJ0 = 1P TT = 10p )

.ENDS LM7815

* Pinouts are the same as 7805.

.SUBCKT LM7818  1    2    3
QT6          23  10  2   Q_NPN 0.1
QT7          5   4   10  Q_NPN 0.1
QT5          7   6   5   Q_NPN 0.1
QT1          1   9   8   Q_NPN 0.1
QT3          11  8   7   Q_NPN 0.1
QT2          11  13  12  Q_NPN 0.1
QT17         1   15  14  Q_NPN 10
C2           10  23      4P
R16          12  5       500
R12          16  2       12.1K
QT18         17  23  16  Q_NPN 0.1
D1           18  19  	 D_D 
R11          20  21      850
R5           22  3       100
QT14         24  18  2   Q_NPN 0.1
R21          6   2       2.67K
R20          3   6       9.142K
DZ2          25  26      D_5V1 
R19          1   26      16K
R18          14  3       250M
R17          25  14      380
R15          25  15      1.62K
QT16         1   20  15  Q_NPN 1
QT15         2   24  21  Q_PNP 0.1 
*OFF
R14          21  24      4K
C1           27  24      20P
R13          19  2       4K
QT13         24  27  18  Q_NPN 0.1
QT12         20  25  22  Q_NPN 1 
*OFF
QT11         20  28  2   Q_NPN 0.1
*OFF
QT10         20  11  1   Q_PNP 0.1
R10          17  27      16.5K
R9           5   4       1.9K
R8           4   23      26
R7           10  2       1.2K
R6           29  2       1K
QT9          11  11  1   Q_PNP 0.1
QT8          27  16  29  Q_NPN 0.1
QT4          15  6   17  Q_NPN 0.1
DZ1          2   9       D_5V6
R4           1   9       80K
R3           28  2       830
R2           13  28      4.97K
R1           8   13      7K

.MODEL D_5V1 D( IS=10F N=1.16 BV=5.1 IBV=0.5M CJ0 = 1P TT = 10p )
.MODEL D_5V6 D( IS=10F N=1.16 BV=5.6 IBV=5U CJ0 = 1P TT = 10p )
.MODEL Q_NPN NPN( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+       TF=10P TR=1N )
.MODEL Q_PNP PNP( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+      TF=10P TR=1N )
.MODEL D_D D( IS=1F N=1.16 CJ0 = 1P TT = 10p )

.ENDS LM7818

* Pinouts are the same as 7805.

.SUBCKT LM7824  1    2    3
QT6          23  10  2   Q_NPN 0.1
QT7          5   4   10  Q_NPN 0.1
QT5          7   6   5   Q_NPN 0.1
QT1          1   9   8   Q_NPN 0.1
QT3          11  8   7   Q_NPN 0.1
QT2          11  13  12  Q_NPN 0.1
QT17         1   15  14  Q_NPN 10
C2           10  23      4P
R16          12  5       500
R12          16  2       12.1K
QT18         17  23  16  Q_NPN 0.1
D1           18  19  	 D_D 
R11          20  21      850
R5           22  3       100
QT14         24  18  2   Q_NPN 0.1
R21          6   2       2.67K
R20          3   6       13.07K
DZ2          25  26      D_5V1 
R19          1   26      16K
R18          14  3       250M
R17          25  14      380
R15          25  15      1.62K
QT16         1   20  15  Q_NPN 1
QT15         2   24  21  Q_PNP 0.1 
*OFF
R14          21  24      4K
C1           27  24      20P
R13          19  2       4K
QT13         24  27  18  Q_NPN 0.1
QT12         20  25  22  Q_NPN 1 
*OFF
QT11         20  28  2   Q_NPN 0.1
*OFF
QT10         20  11  1   Q_PNP 0.1
R10          17  27      16.5K
R9           5   4       1.9K
R8           4   23      26
R7           10  2       1.2K
R6           29  2       1K
QT9          11  11  1   Q_PNP 0.1
QT8          27  16  29  Q_NPN 0.1
QT4          15  6   17  Q_NPN 0.1
DZ1          2   9       D_5V6
R4           1   9       80K
R3           28  2       830
R2           13  28      4.97K
R1           8   13      7K

.MODEL D_5V1 D( IS=10F N=1.16 BV=5.1 IBV=0.5M CJ0 = 1P TT = 10p )
.MODEL D_5V6 D( IS=10F N=1.16 BV=5.6 IBV=5U CJ0 = 1P TT = 10p )
.MODEL Q_NPN NPN( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+       TF=10P TR=1N )
.MODEL Q_PNP PNP( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+      TF=10P TR=1N )
.MODEL D_D D( IS=1F N=1.16 CJ0 = 1P TT = 10p )

.ENDS LM7824


* Identical.

.SUBCKT LM7905  1    2    3            

DD4           4   5   D_6V3_0 
DD2           6   2   D_3V9_0 
DD1           7   2   D_4V7_0 
DD3           8   3   D_6V3_0 
C2            9  10  5P
C1            2   9  15P
QTU15         10   9   3   Q_PNP_0 1.000
R17          11  12  4.2K
QTU22          3  10  13   Q_NPN_0 3.000
R18           8   5  15.65K
R20          13  14  1K
R19           4  14  75
QTU31         12  11   4   Q_NPN_1 1.000
R16          15   1  160
R24          16   1  1.8k
C3           17   1  10P
QTU30         18  12  15   Q_NPN_1 1.000
QTU29         10  16   1   Q_NPN_1 1.000
R15          19   1  400
QTU28         10  20  19   Q_NPN_1 1.000
R14          21   1  200
QTU27         17  20  21   Q_NPN_1 1.000
R11          22  23  1K
R10          24  25  1K
QTU19         18  27  26   Q_NPN_1 1.000
R9            2  18  7.1K
QTU8          16  18   2   Q_PNP_0 1.000
QTU7          28  18   2   Q_PNP_0 1.000
QTU6          18  18   2   Q_PNP_0 1.000
QTU5          11  29   2   Q_PNP_0 1.000
QTU4          20  29   2   Q_PNP_0 1.000
QTU3           1  29   2   Q_PNP_0 1.000
QTU2           1  29   2   Q_PNP_0 1.000
R13          28   1  400
R12          30   1  400
QTU18         29  29  31   Q_NPN_1 1.000
QTU1          29  29   2   Q_PNP_0 1.000
R6           31  32  6.5K
R7           32  27  5.6K
R8           27  26  950
QTU10         33   6  26   Q_PNP_0 1.000
QTU17         34  35  33   Q_PNP_0 1.000
R5           36   1  2K
QTU24         34  34  36   Q_NPN_1 1.000
R1           37   6  6.3K
R2           37  38  670
R3           38  35  550
QTU9          38  35   6   Q_PNP_0 1.000
R4           39   1  2K
QTU23         35  34  39   Q_NPN_1 1.000
QTU16          1   7  35   Q_PNP_0 1.000
JT1           7   1   1  J_2N3458_N 
QTU14          3  17  23   Q_PNP_0 1.000
QTU13         17  17  23   Q_PNP_0 1.000
QTU12         17  17  25   Q_PNP_0 1.000
QTU11          9  17  25   Q_PNP_0 1.000
QTU32          3  13  14   Q_NPN_2 10.000
QTU26          9  20  28   Q_NPN_1 1.000
QTU25         20  20  30   Q_NPN_1 1.000
QTU21          2  40  22   Q_NPN_1 1.000
QTU20          2  37  24   Q_NPN_1 1.000
R21           2  40  4.29K
R22          40   3  500
R23          14   1  500M

.MODEL J_2N3458_N NJF( VTO=-3.05 BETA=699.53U LAMBDA=6M RD=1 RS=1 
+      CGD=2.81P CGS=2.91P M=227.1M PB=500M IS=114.41F 
+      VTOTC=-2.5M BETATCE=-500M KF=0 AF=1 )
.MODEL D_6V3_0  D( IS=10F N=1.24 BV=6.3 IBV=1M CJ0 = 1P TT = 10p )
.MODEL D_3V9_0  D( IS=10F N=1.24 BV=3.9 IBV=1M CJ0 = 1P TT = 10p )
.MODEL D_4V7_0  D( IS=10F N=1.24 BV=4.7 IBV=1M CJ0 = 1P TT = 10p )
.MODEL Q_PNP_0  PNP( IS=10F NF=1.04 NR=1.04 BF=50 CJC=1P CJE=2P
+      TF=10P TR=1N VAF=45)
.MODEL Q_NPN_0  NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.MODEL Q_NPN_1  NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.MODEL Q_NPN_2  NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.ENDS LM7905

* Identical.

.SUBCKT LM7906  1    2    3            

DD4           4   5   D_6V3_0 
DD2           6   2   D_3V9_0 
DD1           7   2   D_4V7_0 
DD3           8   3   D_6V3_0 
C2            9  10  5P
C1            2   9  15P
QTU15         10   9   3   Q_PNP_0 1.000
R17          11  12  4.2K
QTU22          3  10  13   Q_NPN_0 3.000
R18           8   5  15.65K
R20          13  14  1K
R19           4  14  75
QTU31         12  11   4   Q_NPN_1 1.000
R16          15   1  160
R24          16   1  1.8k
C3           17   1  10P
QTU30         18  12  15   Q_NPN_1 1.000
QTU29         10  16   1   Q_NPN_1 1.000
R15          19   1  400
QTU28         10  20  19   Q_NPN_1 1.000
R14          21   1  200
QTU27         17  20  21   Q_NPN_1 1.000
R11          22  23  1K
R10          24  25  1K
QTU19         18  27  26   Q_NPN_1 1.000
R9            2  18  7.1K
QTU8          16  18   2   Q_PNP_0 1.000
QTU7          28  18   2   Q_PNP_0 1.000
QTU6          18  18   2   Q_PNP_0 1.000
QTU5          11  29   2   Q_PNP_0 1.000
QTU4          20  29   2   Q_PNP_0 1.000
QTU3           1  29   2   Q_PNP_0 1.000
QTU2           1  29   2   Q_PNP_0 1.000
R13          28   1  400
R12          30   1  400
QTU18         29  29  31   Q_NPN_1 1.000
QTU1          29  29   2   Q_PNP_0 1.000
R6           31  32  6.5K
R7           32  27  5.6K
R8           27  26  950
QTU10         33   6  26   Q_PNP_0 1.000
QTU17         34  35  33   Q_PNP_0 1.000
R5           36   1  2K
QTU24         34  34  36   Q_NPN_1 1.000
R1           37   6  6.3K
R2           37  38  670
R3           38  35  550
QTU9          38  35   6   Q_PNP_0 1.000
R4           39   1  2K
QTU23         35  34  39   Q_NPN_1 1.000
QTU16          1   7  35   Q_PNP_0 1.000
JT1           7   1   1  J_2N3458_N 
QTU14          3  17  23   Q_PNP_0 1.000
QTU13         17  17  23   Q_PNP_0 1.000
QTU12         17  17  25   Q_PNP_0 1.000
QTU11          9  17  25   Q_PNP_0 1.000
QTU32          3  13  14   Q_NPN_2 10.000
QTU26          9  20  28   Q_NPN_1 1.000
QTU25         20  20  30   Q_NPN_1 1.000
QTU21          2  40  22   Q_NPN_1 1.000
QTU20          2  37  24   Q_NPN_1 1.000
R21           2  40  4.29K
R22          40   3  1.17K
R23          14   1  500M

.MODEL J_2N3458_N NJF( VTO=-3.05 BETA=699.53U LAMBDA=6M RD=1 RS=1 
+      CGD=2.81P CGS=2.91P M=227.1M PB=500M IS=114.41F 
+      VTOTC=-2.5M BETATCE=-500M KF=0 AF=1 )
.MODEL D_6V3_0  D( IS=10F N=1.24 BV=6.3 IBV=1M CJ0 = 1P TT = 10p )
.MODEL D_3V9_0  D( IS=10F N=1.24 BV=3.9 IBV=1M CJ0 = 1P TT = 10p )
.MODEL D_4V7_0  D( IS=10F N=1.24 BV=4.7 IBV=1M CJ0 = 1P TT = 10p )
.MODEL Q_PNP_0  PNP( IS=10F NF=1.04 NR=1.04 BF=50 CJC=1P CJE=2P
+      TF=10P TR=1N VAF=45)
.MODEL Q_NPN_0  NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.MODEL Q_NPN_1  NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.MODEL Q_NPN_2  NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.ENDS LM7906

* Identical.

.SUBCKT LM7908  1    2    3            

DD4           4   5   D_6V3_0 
DD2           6   2   D_3V9_0 
DD1           7   2   D_4V7_0 
DD3           8   3   D_6V3_0 
C2            9  10  5P
C1            2   9  15P
QTU15         10   9   3   Q_PNP_0 1.000
R17          11  12  4.2K
QTU22          3  10  13   Q_NPN_0 3.000
R18           8   5  15.65K
R20          13  14  1K
R19           4  14  75
QTU31         12  11   4   Q_NPN_1 1.000
R16          15   1  160
R24          16   1  1.8k
C3           17   1  10P
QTU30         18  12  15   Q_NPN_1 1.000
QTU29         10  16   1   Q_NPN_1 1.000
R15          19   1  400
QTU28         10  20  19   Q_NPN_1 1.000
R14          21   1  200
QTU27         17  20  21   Q_NPN_1 1.000
R11          22  23  1K
R10          24  25  1K
QTU19         18  27  26   Q_NPN_1 1.000
R9            2  18  7.1K
QTU8          16  18   2   Q_PNP_0 1.000
QTU7          28  18   2   Q_PNP_0 1.000
QTU6          18  18   2   Q_PNP_0 1.000
QTU5          11  29   2   Q_PNP_0 1.000
QTU4          20  29   2   Q_PNP_0 1.000
QTU3           1  29   2   Q_PNP_0 1.000
QTU2           1  29   2   Q_PNP_0 1.000
R13          28   1  400
R12          30   1  400
QTU18         29  29  31   Q_NPN_1 1.000
QTU1          29  29   2   Q_PNP_0 1.000
R6           31  32  6.5K
R7           32  27  5.6K
R8           27  26  950
QTU10         33   6  26   Q_PNP_0 1.000
QTU17         34  35  33   Q_PNP_0 1.000
R5           36   1  2K
QTU24         34  34  36   Q_NPN_1 1.000
R1           37   6  6.3K
R2           37  38  670
R3           38  35  550
QTU9          38  35   6   Q_PNP_0 1.000
R4           39   1  2K
QTU23         35  34  39   Q_NPN_1 1.000
QTU16          1   7  35   Q_PNP_0 1.000
JT1           7   1   1  J_2N3458_N 
QTU14          3  17  23   Q_PNP_0 1.000
QTU13         17  17  23   Q_PNP_0 1.000
QTU12         17  17  25   Q_PNP_0 1.000
QTU11          9  17  25   Q_PNP_0 1.000
QTU32          3  13  14   Q_NPN_2 10.000
QTU26          9  20  28   Q_NPN_1 1.000
QTU25         20  20  30   Q_NPN_1 1.000
QTU21          2  40  22   Q_NPN_1 1.000
QTU20          2  37  24   Q_NPN_1 1.000
R21           2  40  4.29K
R22          40   3  3.28K
R23          14   1  500M

.MODEL J_2N3458_N NJF( VTO=-3.05 BETA=699.53U LAMBDA=6M RD=1 RS=1 
+      CGD=2.81P CGS=2.91P M=227.1M PB=500M IS=114.41F 
+      VTOTC=-2.5M BETATCE=-500M KF=0 AF=1 )
.MODEL D_6V3_0  D( IS=10F N=1.24 BV=6.3 IBV=1M CJ0 = 1P TT = 10p )
.MODEL D_3V9_0  D( IS=10F N=1.24 BV=3.9 IBV=1M CJ0 = 1P TT = 10p )
.MODEL D_4V7_0  D( IS=10F N=1.24 BV=4.7 IBV=1M CJ0 = 1P TT = 10p )
.MODEL Q_PNP_0  PNP( IS=10F NF=1.04 NR=1.04 BF=50 CJC=1P CJE=2P
+      TF=10P TR=1N VAF=45)
.MODEL Q_NPN_0  NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.MODEL Q_NPN_1  NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.MODEL Q_NPN_2  NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.ENDS LM7908

* Identical.

.SUBCKT LM7909  1    2    3            

DD4           4   5   D_6V3_0 
DD2           6   2   D_3V9_0 
DD1           7   2   D_4V7_0 
DD3           8   3   D_6V3_0 
C2            9  10  5P
C1            2   9  15P
QTU15         10   9   3   Q_PNP_0 1.000
R17          11  12  4.2K
QTU22          3  10  13   Q_NPN_0 3.000
R18           8   5  15.65K
R20          13  14  1K
R19           4  14  75
QTU31         12  11   4   Q_NPN_1 1.000
R16          15   1  160
R24          16   1  1.8k
C3           17   1  10P
QTU30         18  12  15   Q_NPN_1 1.000
QTU29         10  16   1   Q_NPN_1 1.000
R15          19   1  400
QTU28         10  20  19   Q_NPN_1 1.000
R14          21   1  200
QTU27         17  20  21   Q_NPN_1 1.000
R11          22  23  1K
R10          24  25  1K
QTU19         18  27  26   Q_NPN_1 1.000
R9            2  18  7.1K
QTU8          16  18   2   Q_PNP_0 1.000
QTU7          28  18   2   Q_PNP_0 1.000
QTU6          18  18   2   Q_PNP_0 1.000
QTU5          11  29   2   Q_PNP_0 1.000
QTU4          20  29   2   Q_PNP_0 1.000
QTU3           1  29   2   Q_PNP_0 1.000
QTU2           1  29   2   Q_PNP_0 1.000
R13          28   1  400
R12          30   1  400
QTU18         29  29  31   Q_NPN_1 1.000
QTU1          29  29   2   Q_PNP_0 1.000
R6           31  32  6.5K
R7           32  27  5.6K
R8           27  26  950
QTU10         33   6  26   Q_PNP_0 1.000
QTU17         34  35  33   Q_PNP_0 1.000
R5           36   1  2K
QTU24         34  34  36   Q_NPN_1 1.000
R1           37   6  6.3K
R2           37  38  670
R3           38  35  550
QTU9          38  35   6   Q_PNP_0 1.000
R4           39   1  2K
QTU23         35  34  39   Q_NPN_1 1.000
QTU16          1   7  35   Q_PNP_0 1.000
JT1           7   1   1  J_2N3458_N 
QTU14          3  17  23   Q_PNP_0 1.000
QTU13         17  17  23   Q_PNP_0 1.000
QTU12         17  17  25   Q_PNP_0 1.000
QTU11          9  17  25   Q_PNP_0 1.000
QTU32          3  13  14   Q_NPN_2 10.000
QTU26          9  20  28   Q_NPN_1 1.000
QTU25         20  20  30   Q_NPN_1 1.000
QTU21          2  40  22   Q_NPN_1 1.000
QTU20          2  37  24   Q_NPN_1 1.000
R21           2  40  4.29K
R22          40   3  4.33K
R23          14   1  500M

.MODEL J_2N3458_N NJF( VTO=-3.05 BETA=699.53U LAMBDA=6M RD=1 RS=1 
+      CGD=2.81P CGS=2.91P M=227.1M PB=500M IS=114.41F 
+      VTOTC=-2.5M BETATCE=-500M KF=0 AF=1 )
.MODEL D_6V3_0  D( IS=10F N=1.24 BV=6.3 IBV=1M CJ0 = 1P TT = 10p )
.MODEL D_3V9_0  D( IS=10F N=1.24 BV=3.9 IBV=1M CJ0 = 1P TT = 10p )
.MODEL D_4V7_0  D( IS=10F N=1.24 BV=4.7 IBV=1M CJ0 = 1P TT = 10p )
.MODEL Q_PNP_0  PNP( IS=10F NF=1.04 NR=1.04 BF=50 CJC=1P CJE=2P
+      TF=10P TR=1N VAF=45)
.MODEL Q_NPN_0  NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.MODEL Q_NPN_1  NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.MODEL Q_NPN_2  NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.ENDS LM7909

* Identical.

.SUBCKT LM79XX Input Output Ground PARAMS:
+       Av_feedback=1660, R1_Value=4615,
+       Rbg_Tc1=8.13E-5, Rbg_Tc2=0.0,
+       Rout_Value=0.01, Rreg_Value=9.1k ;1.2k
*
* SERIES 3-TERMINAL NEGATIVE REGULATOR
*
* Note: This regulator is based on the LM79XX series of
*       regulators (also the LM120 and LM320).  The
*       LM79XX regulators are unstable and will
*       oscillate unless a 1 uFarad solid tantalum
*       capacitor is placed on the output with an ESR
*       betweed .5 and 1.5.  This model is stable without
*       a capacitor on the output.  When performing
*       simulations a 1 uFarad capacitor should still be
*       placed on the output.  However, it it not necessary
*       to include a resistor in series with this capacitor
*       to model the ESR of the capacitor.  See the
*       comments and circuit description of the x_LM78XX
*       regulator for more information on this model.
*
* Band-gap voltage source:
*
Vbg 100 0 DC -7.4V
Sbg 100 101 Ground Input  Sbg1
Rbg 101 0 Rbg1 1
.MODEL Rbg1 RES (Tc1={Rbg_Tc1},Tc2={Rbg_Tc2})
Ebg 102 0 Input Ground  1
Rreg 102 101 {Rreg_Value}
.MODEL Sbg1 VSWITCH (Ron=1 Roff=1MEG Von=3.7 Voff=3)
*
* Feedback stage
*
Rfb 9 8 1MEG
Cfb 8 Ground 265PF
* Eopamp 105 0 VALUE={2250*v(101,0)+Av_feedback*v(Ground,8)}
Vgainf 200 0 {Av_feedback}
Rgainf 200 0 1
Eopamp 105 0 POLY(3),(101,0),(Ground,8),(200,0) 0 2250 0 0 0 0 0 0 1
Ro 105 106 1k
D1 108 106 Dlim
D2 106 107 Dlim
.MODEL Dlim D (Vj=0.7)
Vl1 108 102 DC 1
Vl2 0 107 DC 1
*
* Quiescent current modelling
*
Gq (Ground,Input),(9,Input) 9.0E-7
R1 9 Ground {R1_Value} TC=0.001
Fl (Ground,0) Vmon 3.0E-4
*
* Output Stage
*
Q1 9 5 6 Npn1
Q2 9 6 7 Npn1 10
.MODEL Npn1 NPN (Bf=50 Is=1E-14)
* Efb 4 Ground VALUE={v(Input,Ground)+v(0,106)}
Efb 4 Ground POLY(2)  (Input,Ground) (0,106) 0 1 1
Rb 4 5 1k TC=0.003
Re 6 7 2k
Rsc 7 Input 0.13 TC=1.136E-3,-7.806E-6
Rout 9 Imon {Rout_Value}
Vmon Imon Output DC 0.0
*
* Current Limit
*
Qcl1 54 52 53 Npn1
Qcl3 Input 54 5 Pnp1
.MODEL Pnp1 PNP (Bf=250 Is=1E-14)
Rcl3 5 54 1.8k
Qcl2 52 52 51 Npn1
Veset 53 Input DC 0.3v
Ibias Input 52 DC 300u
Rcl1 50 51 20k
Rcl2 51 7 115
Dz1 50 9 Dz
.MODEL Dz D (Is=0.05p Rs=3 Bv=7.11 Ibv=0.05u)
.ENDS


.SUBCKT LM7912  INPUT  GROUND OUTPUT
x1 Input Output Ground  LM79XX PARAMS:
+     Av_feedback=694, R1_Value=11076,
+     Rbg_Tc1=-9.50E-7, Rbg_Tc2=-6.53E-7,
+     Rout_Value=0.01, Rreg_Value=9.1k
.ENDS



* Identical.

.SUBCKT LM7915  1    2    3            

DD4           4   5   D_6V3_0 
DD2           6   2   D_3V9_0 
DD1           7   2   D_4V7_0 
DD3           8   3   D_6V3_0 
C2            9  10  5P
C1            2   9  15P
QTU15         10   9   3   Q_PNP_0 1.000
R17          11  12  4.2K
QTU22          3  10  13   Q_NPN_0 3.000
R18           8   5  15.65K
R20          13  14  1K
R19           4  14  75
QTU31         12  11   4   Q_NPN_1 1.000
R16          15   1  160
R24          16   1  1.8k
C3           17   1  10P
QTU30         18  12  15   Q_NPN_1 1.000
QTU29         10  16   1   Q_NPN_1 1.000
R15          19   1  400
QTU28         10  20  19   Q_NPN_1 1.000
R14          21   1  200
QTU27         17  20  21   Q_NPN_1 1.000
R11          22  23  1K
R10          24  25  1K
QTU19         18  27  26   Q_NPN_1 1.000
R9            2  18  7.1K
QTU8          16  18   2   Q_PNP_0 1.000
QTU7          28  18   2   Q_PNP_0 1.000
QTU6          18  18   2   Q_PNP_0 1.000
QTU5          11  29   2   Q_PNP_0 1.000
QTU4          20  29   2   Q_PNP_0 1.000
QTU3           1  29   2   Q_PNP_0 1.000
QTU2           1  29   2   Q_PNP_0 1.000
R13          28   1  400
R12          30   1  400
QTU18         29  29  31   Q_NPN_1 1.000
QTU1          29  29   2   Q_PNP_0 1.000
R6           31  32  6.5K
R7           32  27  5.6K
R8           27  26  950
QTU10         33   6  26   Q_PNP_0 1.000
QTU17         34  35  33   Q_PNP_0 1.000
R5           36   1  2K
QTU24         34  34  36   Q_NPN_1 1.000
R1           37   6  6.3K
R2           37  38  670
R3           38  35  550
QTU9          38  35   6   Q_PNP_0 1.000
R4           39   1  2K
QTU23         35  34  39   Q_NPN_1 1.000
QTU16          1   7  35   Q_PNP_0 1.000
JT1           7   1   1  J_2N3458_N 
QTU14          3  17  23   Q_PNP_0 1.000
QTU13         17  17  23   Q_PNP_0 1.000
QTU12         17  17  25   Q_PNP_0 1.000
QTU11          9  17  25   Q_PNP_0 1.000
QTU32          3  13  14   Q_NPN_2 10.000
QTU26          9  20  28   Q_NPN_1 1.000
QTU25         20  20  30   Q_NPN_1 1.000
QTU21          2  40  22   Q_NPN_1 1.000
QTU20          2  37  24   Q_NPN_1 1.000
R21           2  40  4.29K
R22          40   3  10.66K
R23          14   1  500M

.MODEL J_2N3458_N NJF( VTO=-3.05 BETA=699.53U LAMBDA=6M RD=1 RS=1 
+      CGD=2.81P CGS=2.91P M=227.1M PB=500M IS=114.41F 
+      VTOTC=-2.5M BETATCE=-500M KF=0 AF=1 )
.MODEL D_6V3_0  D( IS=10F N=1.24 BV=6.3 IBV=1M CJ0 = 1P TT = 10p )
.MODEL D_3V9_0  D( IS=10F N=1.24 BV=3.9 IBV=1M CJ0 = 1P TT = 10p )
.MODEL D_4V7_0  D( IS=10F N=1.24 BV=4.7 IBV=1M CJ0 = 1P TT = 10p )
.MODEL Q_PNP_0  PNP( IS=10F NF=1.04 NR=1.04 BF=50 CJC=1P CJE=2P
+      TF=10P TR=1N VAF=45)
.MODEL Q_NPN_0  NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.MODEL Q_NPN_1  NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.MODEL Q_NPN_2  NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.ENDS LM7915

* Identical but PIN 2 is now ADJUST instead of GND.
* LM117 seems to be the same model.

* Identical.

.SUBCKT LM7918  1    2    3            

DD4           4   5   D_6V3_0 
DD2           6   2   D_3V9_0 
DD1           7   2   D_4V7_0 
DD3           8   3   D_6V3_0 
C2            9  10  5P
C1            2   9  15P
QTU15         10   9   3   Q_PNP_0 1.000
R17          11  12  4.2K
QTU22          3  10  13   Q_NPN_0 3.000
R18           8   5  15.65K
R20          13  14  1K
R19           4  14  75
QTU31         12  11   4   Q_NPN_1 1.000
R16          15   1  160
R24          16   1  1.8k
C3           17   1  10P
QTU30         18  12  15   Q_NPN_1 1.000
QTU29         10  16   1   Q_NPN_1 1.000
R15          19   1  400
QTU28         10  20  19   Q_NPN_1 1.000
R14          21   1  200
QTU27         17  20  21   Q_NPN_1 1.000
R11          22  23  1K
R10          24  25  1K
QTU19         18  27  26   Q_NPN_1 1.000
R9            2  18  7.1K
QTU8          16  18   2   Q_PNP_0 1.000
QTU7          28  18   2   Q_PNP_0 1.000
QTU6          18  18   2   Q_PNP_0 1.000
QTU5          11  29   2   Q_PNP_0 1.000
QTU4          20  29   2   Q_PNP_0 1.000
QTU3           1  29   2   Q_PNP_0 1.000
QTU2           1  29   2   Q_PNP_0 1.000
R13          28   1  400
R12          30   1  400
QTU18         29  29  31   Q_NPN_1 1.000
QTU1          29  29   2   Q_PNP_0 1.000
R6           31  32  6.5K
R7           32  27  5.6K
R8           27  26  950
QTU10         33   6  26   Q_PNP_0 1.000
QTU17         34  35  33   Q_PNP_0 1.000
R5           36   1  2K
QTU24         34  34  36   Q_NPN_1 1.000
R1           37   6  6.3K
R2           37  38  670
R3           38  35  550
QTU9          38  35   6   Q_PNP_0 1.000
R4           39   1  2K
QTU23         35  34  39   Q_NPN_1 1.000
QTU16          1   7  35   Q_PNP_0 1.000
JT1           7   1   1  J_2N3458_N 
QTU14          3  17  23   Q_PNP_0 1.000
QTU13         17  17  23   Q_PNP_0 1.000
QTU12         17  17  25   Q_PNP_0 1.000
QTU11          9  17  25   Q_PNP_0 1.000
QTU32          3  13  14   Q_NPN_2 10.000
QTU26          9  20  28   Q_NPN_1 1.000
QTU25         20  20  30   Q_NPN_1 1.000
QTU21          2  40  22   Q_NPN_1 1.000
QTU20          2  37  24   Q_NPN_1 1.000
R21           2  40  4.29K
R22          40   3  13.83K
R23          14   1  500M

.MODEL J_2N3458_N NJF( VTO=-3.05 BETA=699.53U LAMBDA=6M RD=1 RS=1 
+      CGD=2.81P CGS=2.91P M=227.1M PB=500M IS=114.41F 
+      VTOTC=-2.5M BETATCE=-500M KF=0 AF=1 )
.MODEL D_6V3_0  D( IS=10F N=1.24 BV=6.3 IBV=1M CJ0 = 1P TT = 10p )
.MODEL D_3V9_0  D( IS=10F N=1.24 BV=3.9 IBV=1M CJ0 = 1P TT = 10p )
.MODEL D_4V7_0  D( IS=10F N=1.24 BV=4.7 IBV=1M CJ0 = 1P TT = 10p )
.MODEL Q_PNP_0  PNP( IS=10F NF=1.04 NR=1.04 BF=50 CJC=1P CJE=2P
+      TF=10P TR=1N VAF=45)
.MODEL Q_NPN_0  NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.MODEL Q_NPN_1  NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.MODEL Q_NPN_2  NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.ENDS LM7918

* Identical.

.SUBCKT LM7924  1    2    3            

DD4           4   5   D_6V3_0 
DD2           6   2   D_3V9_0 
DD1           7   2   D_4V7_0 
DD3           8   3   D_6V3_0 
C2            9  10  5P
C1            2   9  15P
QTU15         10   9   3   Q_PNP_0 1.000
R17          11  12  4.2K
QTU22          3  10  13   Q_NPN_0 3.000
R18           8   5  15.65K
R20          13  14  1K
R19           4  14  75
QTU31         12  11   4   Q_NPN_1 1.000
R16          15   1  160
R24          16   1  1.8k
C3           17   1  10P
QTU30         18  12  15   Q_NPN_1 1.000
QTU29         10  16   1   Q_NPN_1 1.000
R15          19   1  400
QTU28         10  20  19   Q_NPN_1 1.000
R14          21   1  200
QTU27         17  20  21   Q_NPN_1 1.000
R11          22  23  1K
R10          24  25  1K
QTU19         18  27  26   Q_NPN_1 1.000
R9            2  18  7.1K
QTU8          16  18   2   Q_PNP_0 1.000
QTU7          28  18   2   Q_PNP_0 1.000
QTU6          18  18   2   Q_PNP_0 1.000
QTU5          11  29   2   Q_PNP_0 1.000
QTU4          20  29   2   Q_PNP_0 1.000
QTU3           1  29   2   Q_PNP_0 1.000
QTU2           1  29   2   Q_PNP_0 1.000
R13          28   1  400
R12          30   1  400
QTU18         29  29  31   Q_NPN_1 1.000
QTU1          29  29   2   Q_PNP_0 1.000
R6           31  32  6.5K
R7           32  27  5.6K
R8           27  26  950
QTU10         33   6  26   Q_PNP_0 1.000
QTU17         34  35  33   Q_PNP_0 1.000
R5           36   1  2K
QTU24         34  34  36   Q_NPN_1 1.000
R1           37   6  6.3K
R2           37  38  670
R3           38  35  550
QTU9          38  35   6   Q_PNP_0 1.000
R4           39   1  2K
QTU23         35  34  39   Q_NPN_1 1.000
QTU16          1   7  35   Q_PNP_0 1.000
JT1           7   1   1  J_2N3458_N 
QTU14          3  17  23   Q_PNP_0 1.000
QTU13         17  17  23   Q_PNP_0 1.000
QTU12         17  17  25   Q_PNP_0 1.000
QTU11          9  17  25   Q_PNP_0 1.000
QTU32          3  13  14   Q_NPN_2 10.000
QTU26          9  20  28   Q_NPN_1 1.000
QTU25         20  20  30   Q_NPN_1 1.000
QTU21          2  40  22   Q_NPN_1 1.000
QTU20          2  37  24   Q_NPN_1 1.000
R21           2  40  4.29K
R22          40   3  20.16K
R23          14   1  500M

.MODEL J_2N3458_N NJF( VTO=-3.05 BETA=699.53U LAMBDA=6M RD=1 RS=1 
+      CGD=2.81P CGS=2.91P M=227.1M PB=500M IS=114.41F 
+      VTOTC=-2.5M BETATCE=-500M KF=0 AF=1 )
.MODEL D_6V3_0  D( IS=10F N=1.24 BV=6.3 IBV=1M CJ0 = 1P TT = 10p )
.MODEL D_3V9_0  D( IS=10F N=1.24 BV=3.9 IBV=1M CJ0 = 1P TT = 10p )
.MODEL D_4V7_0  D( IS=10F N=1.24 BV=4.7 IBV=1M CJ0 = 1P TT = 10p )
.MODEL Q_PNP_0  PNP( IS=10F NF=1.04 NR=1.04 BF=50 CJC=1P CJE=2P
+      TF=10P TR=1N VAF=45)
.MODEL Q_NPN_0  NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.MODEL Q_NPN_1  NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.MODEL Q_NPN_2  NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.ENDS LM7924

.SUBCKT LM317    1    2    3
D4            4   3  D_Z6V0
D3            5   6  D_Z6V3
D2            7   1  D_Z6V3
D1            3   8  D_Z6V3
QT26          1  10   9  Q_NPN 20.0
QT25          1  11  10  Q_NPN 2.0
QT24_2       13  12   5  Q_NPN 0.1
QT24         13  12  14  Q_NPN 0.1
QT23         17  16  15  Q_NPN 1.0
QT21         19  18   3  Q_NPN 0.1
QT19         21   3  20  Q_NPN 1.0
QT17         23   3  22  Q_NPN 0.1
QT13          1  25  24  Q_NPN 0.1
QT11         16  27  26  Q_NPN 0.1
QT7          30  29  28  Q_NPN 0.1
QT5          29  31   3  Q_NPN 0.1
QT3          33  31  32  Q_NPN 0.1
QT22_2       17  17   1  Q_PNP 1.0
QT22         16  17   1  Q_PNP 1.0
QT20          3  19  16  Q_PNP 0.1
QT18         21  21  16  Q_PNP 0.1
QT16         23  21  16  Q_PNP 0.1
QT15          3  23  25  Q_PNP 0.1
QT12          3  24  16  Q_PNP 0.1
QT9          27  30  34  Q_PNP 0.1
QT6           3  29  34  Q_PNP 0.1
QT14         25  33  35  Q_PNP 0.1
QT10         16  33  36  Q_PNP 0.1
QT8          34  33  37  Q_PNP 0.1
QT4          31  33  38  Q_PNP 0.1
QT2          33  33  39  Q_PNP 0.1
R27           4   2  50
R26           9   3  100M
R25           9  14  2
R24           5  14  160
R23           7   6  18K
R22          10   3  160
R21          12  13  400
R20          18  13  13K
R19          16  11  370
R18          15  10  130
R17          16  12  12K
C3           19  18  5P
R16          16  19  6.7K
R15          20  22  2.4K
R14          22   4  12K
C2           23   4  30P
C1           23   3  30P
R13          24   3  5.1K
R12          26   3  72
R11          27   3  5.8K
R10          28   3  4.1K
R9           32   3  180
R8           34  30  12.4K
R7           31  29  130
R6            8  31  100K
R5            1  35  5.6K
R4            1  36  82
R3            1  37  190
R2            1  38  310
R1            1  39  310
JT1           1   3   8  J_N

.MODEL D_Z6V0 D( IS=10F N=1.04 BV=6.0 IBV=1M CJ0 = 1P TT = 10p )
.MODEL D_Z6V3 D( IS=10F N=1.04 BV=6.3 IBV=1M CJ0 = 1P TT = 10p )
.MODEL Q_NPN NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.MODEL Q_PNP PNP( IS=10F NF=1.04 NR=1.04 BF=50 CJC=1P CJE=2P
+      TF=10P TR=1N VAF=45)
.MODEL J_N NJF( VTO=-7 )

.ENDS LM117




* LM7805 model. 
* No need to use .inc - I've set the .asy symbol to remove the need for .inc.
* (I used the symbol of LT1084, just replaced the LT1084 by LMxxxx and LTC.LIB by regulators.lib) 

.SUBCKT LM7805-1 1    2    3
* In GND Out
QT6          23  10  2   Q_NPN 0.1
QT7          5   4   10  Q_NPN 0.1
QT5          7   6   5   Q_NPN 0.1
QT1          1   9   8   Q_NPN 0.1
QT3          11  8   7   Q_NPN 0.1
QT2          11  13  12  Q_NPN 0.1
QT17         1   15  14  Q_NPN 10
C2           10  23      4P
R16          12  5       500
R12          16  2       12.1K
QT18         17  23  16  Q_NPN 0.1
D1           18  19      D_D 
R11          20  21      850
R5           22  3       100
QT14         24  18  2   Q_NPN 0.1
R21          6   2       2.67K
R20          3   6       640
DZ2          25  26      D_5V1 
R19          1   26      16K
R18          14  3       250M
R17          25  14      380
R15          25  15      1.62K
QT16         1   20  15  Q_NPN 1
QT15         2   24  21  Q_PNP 0.1
*OFF
R14          21  24      4K
C1           27  24      20P
R13          19  2       4K
QT13         24  27  18  Q_NPN 0.1
QT12         20  25  22  Q_NPN 1 
*OFF
QT11         20  28  2   Q_NPN 0.1
*OFF
QT10         20  11  1   Q_PNP 0.1
R10          17  27      16.5K
R9           5   4       1.9K
R8           4   23      26
R7           10  2       1.2K
R6           29  2       1K
QT9          11  11  1   Q_PNP 0.1
QT8          27  16  29  Q_NPN 0.1
QT4          15  6   17  Q_NPN 0.1
DZ1          2   9       D_5V6
R4           1   9       80K
R3           28  2       830
R2           13  28      4.97K
R1           8   13      7K

.MODEL D_5V1 D( IS=10F N=1.16 BV=5.1 IBV=0.5M CJ0 = 1P TT = 10p )
.MODEL D_5V6 D( IS=10F N=1.16 BV=5.6 IBV=5U CJ0 = 1P TT = 10p )
.MODEL Q_NPN NPN( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+       TF=10P TR=1N )
.MODEL Q_PNP PNP( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+      TF=10P TR=1N )
.MODEL D_D D( IS=1F N=1.16 CJ0 = 1P TT = 10p )

.ENDS LM7805-1

*==================================
*LM7808C National Semiconductor
* Connections: Input
*                |   Gnd
*                |    |   Output
*                |    |    |
.SUBCKT LM7808C  1    2    3
QT6          23  10  2   Q_NPN 0.1
QT7          5   4   10  Q_NPN 0.1
QT5          7   6   5   Q_NPN 0.1
QT1          1   9   8   Q_NPN 0.1
QT3          11  8   7   Q_NPN 0.1
QT2          11  13  12  Q_NPN 0.1
QT17         1   15  14  Q_NPN 10
C2           10  23      4P
R16          12  5       500
R12          16  2       12.1K
QT18         17  23  16  Q_NPN 0.1
D1           18  19  	 D_D 
R11          20  21      850
R5           22  3       100
QT14         24  18  2   Q_NPN 0.1
R21          6   2       2.67K
R20          3   6       2.6K
DZ2          25  26      D_5V1
R19          1   26      16K
R18          14  3       250M
R17          25  14      380
R15          25  15      1.62K
QT16         1   20  15  Q_NPN 1
QT15         2   24  21  Q_PNP 0.1 
*OFF
R14          21  24      4K
C1           27  24      20P
R13          19  2       4K
QT13         24  27  18  Q_NPN 0.1
QT12         20  25  22  Q_NPN 1 
*OFF
QT11         20  28  2   Q_NPN 0.1
*OFF
QT10         20  11  1   Q_PNP 0.1
R10          17  27      16.5K
R9           5   4       1.9K
R8           4   23      26
R7           10  2       1.2K
R6           29  2       1K
QT9          11  11  1   Q_PNP 0.1
QT8          27  16  29  Q_NPN 0.1
QT4          15  6   17  Q_NPN 0.1
DZ1          2   9       D_5V6
R4           1   9       80K
R3           28  2       830
R2           13  28      4.97K
R1           8   13      7K

.MODEL D_5V1 D( IS=10F N=1.16 BV=5.1 IBV=0.5M CJO = 1P TT = 10p )
.MODEL D_5V6 D( IS=10F N=1.16 BV=5.6 IBV=5U CJO = 1P TT = 10p )
.MODEL Q_NPN NPN( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+       TF=10P TR=1N )
.MODEL Q_PNP PNP( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+      TF=10P TR=1N )
.MODEL D_D D( IS=1F N=1.16 CJO = 1P TT = 10p )

.ENDS LM7808C


* Pinouts are the same as 7805.

.SUBCKT LM7812-1  1    2    3
QT6          23  10  2   Q_NPN 0.1
QT7          5   4   10  Q_NPN 0.1
QT5          7   6   5   Q_NPN 0.1
QT1          1   9   8   Q_NPN 0.1
QT3          11  8   7   Q_NPN 0.1
QT2          11  13  12  Q_NPN 0.1
QT17         1   15  14  Q_NPN 10
C2           10  23      4P
R16          12  5       500
R12          16  2       12.1K
QT18         17  23  16  Q_NPN 0.1
D1           18  19      D_D 
R11          20  21      850
R5           22  3       100
QT14         24  18  2   Q_NPN 0.1
R21          6   2       2.67K
R20          3   6       5.22K
DZ2          25  26      D_5V1 
R19          1   26      16K
R18          14  3       250M
R17          25  14      380
R15          25  15      1.62K
QT16         1   20  15  Q_NPN 1
QT15         2   24  21  Q_PNP 0.1 
*OFF
R14          21  24      4K
C1           27  24      20P
R13          19  2       4K
QT13         24  27  18  Q_NPN 0.1
QT12         20  25  22  Q_NPN 1 
*OFF
QT11         20  28  2   Q_NPN 0.1
*OFF
QT10         20  11  1   Q_PNP 0.1
R10          17  27      16.5K
R9           5   4       1.9K
R8           4   23      26
R7           10  2       1.2K
R6           29  2       1K
QT9          11  11  1   Q_PNP 0.1
QT8          27  16  29  Q_NPN 0.1
QT4          15  6   17  Q_NPN 0.1
DZ1          2   9       D_5V6
R4           1   9       80K
R3           28  2       830
R2           13  28      4.97K
R1           8   13      7K

.MODEL D_5V1 D( IS=10F N=1.16 BV=5.1 IBV=0.5M CJ0 = 1P TT = 10p )
.MODEL D_5V6 D( IS=10F N=1.16 BV=5.6 IBV=5U CJ0 = 1P TT = 10p )
.MODEL Q_NPN NPN( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+       TF=10P TR=1N )
.MODEL Q_PNP PNP( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+      TF=10P TR=1N )
.MODEL D_D D( IS=1F N=1.16 CJ0 = 1P TT = 10p )

.ENDS LM7812-1

* Pinouts are the same as '05

.SUBCKT LM7815-1  1    2    3
QT6          23  10  2   Q_NPN 0.1
QT7          5   4   10  Q_NPN 0.1
QT5          7   6   5   Q_NPN 0.1
QT1          1   9   8   Q_NPN 0.1
QT3          11  8   7   Q_NPN 0.1
QT2          11  13  12  Q_NPN 0.1
QT17         1   15  14  Q_NPN 10
C2           10  23      4P
R16          12  5       500
R12          16  2       12.1K
QT18         17  23  16  Q_NPN 0.1
D1           18  19      D_D 
R11          20  21      850
R5           22  3       100
QT14         24  18  2   Q_NPN 0.1
R21          6   2       2.67K
R20          3   6       7.18K
DZ2          25  26      D_5V1 
R19          1   26      16K
R18          14  3       250M
R17          25  14      380
R15          25  15      1.62K
QT16         1   20  15  Q_NPN 1
QT15         2   24  21  Q_PNP 0.1 
*OFF
R14          21  24      4K
C1           27  24      20P
R13          19  2       4K
QT13         24  27  18  Q_NPN 0.1
QT12         20  25  22  Q_NPN 1 
*OFF
QT11         20  28  2   Q_NPN 0.1
*OFF
QT10         20  11  1   Q_PNP 0.1
R10          17  27      16.5K
R9           5   4       1.9K
R8           4   23      26
R7           10  2       1.2K
R6           29  2       1K
QT9          11  11  1   Q_PNP 0.1
QT8          27  16  29  Q_NPN 0.1
QT4          15  6   17  Q_NPN 0.1
DZ1          2   9       D_5V6
R4           1   9       80K
R3           28  2       830
R2           13  28      4.97K
R1           8   13      7K

.MODEL D_5V1 D( IS=10F N=1.16 BV=5.1 IBV=0.5M CJ0 = 1P TT = 10p )
.MODEL D_5V6 D( IS=10F N=1.16 BV=5.6 IBV=5U CJ0 = 1P TT = 10p )
.MODEL Q_NPN NPN( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+       TF=10P TR=1N )
.MODEL Q_PNP PNP( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+      TF=10P TR=1N )
.MODEL D_D D( IS=1F N=1.16 CJ0 = 1P TT = 10p )

.ENDS LM7815-1





*LM7815C National Semiconductor
* Connections: Input
*                |   Gnd
*                |    |   Output
*                |    |    |
.SUBCKT LM7815C  1    2    3
QT6          23  10  2   Q_NPN 0.1
QT7          5   4   10  Q_NPN 0.1
QT5          7   6   5   Q_NPN 0.1
QT1          1   9   8   Q_NPN 0.1
QT3          11  8   7   Q_NPN 0.1
QT2          11  13  12  Q_NPN 0.1
QT17         1   15  14  Q_NPN 10
C2           10  23      4P
R16          12  5       500
R12          16  2       12.1K
QT18         17  23  16  Q_NPN 0.1
D1           18  19  	 D_D 
R11          20  21      850
R5           22  3       100
QT14         24  18  2   Q_NPN 0.1
R21          6   2       2.67K
R20          3   6       7.18K
DZ2          25  26      D_5V1 
R19          1   26      16K
R18          14  3       250M
R17          25  14      380
R15          25  15      1.62K
QT16         1   20  15  Q_NPN 1
QT15         2   24  21  Q_PNP 0.1 
*OFF
R14          21  24      4K
C1           27  24      20P
R13          19  2       4K
QT13         24  27  18  Q_NPN 0.1
QT12         20  25  22  Q_NPN 1 
*OFF
QT11         20  28  2   Q_NPN 0.1
*OFF
QT10         20  11  1   Q_PNP 0.1
R10          17  27      16.5K
R9           5   4       1.9K
R8           4   23      26
R7           10  2       1.2K
R6           29  2       1K
QT9          11  11  1   Q_PNP 0.1
QT8          27  16  29  Q_NPN 0.1
QT4          15  6   17  Q_NPN 0.1
DZ1          2   9       D_5V6
R4           1   9       80K
R3           28  2       830
R2           13  28      4.97K
R1           8   13      7K

.MODEL D_5V1 D( IS=10F N=1.16 BV=5.1 IBV=0.5M CJO = 1P TT = 10p )
.MODEL D_5V6 D( IS=10F N=1.16 BV=5.6 IBV=5U CJO = 1P TT = 10p )
.MODEL Q_NPN NPN( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+       TF=10P TR=1N )
.MODEL Q_PNP PNP( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+      TF=10P TR=1N )
.MODEL D_D D( IS=1F N=1.16 CJO = 1P TT = 10p )

.ENDS LM7815C

*LM7824C National Semiconductor
* Connections: Input
*                |   Gnd
*                |    |   Output
*                |    |    |
.SUBCKT LM7824C  1    2    3
QT6          23  10  2   Q_NPN 0.1
QT7          5   4   10  Q_NPN 0.1
QT5          7   6   5   Q_NPN 0.1
QT1          1   9   8   Q_NPN 0.1
QT3          11  8   7   Q_NPN 0.1
QT2          11  13  12  Q_NPN 0.1
QT17         1   15  14  Q_NPN 10
C2           10  23      4P
R16          12  5       500
R12          16  2       12.1K
QT18         17  23  16  Q_NPN 0.1
D1           18  19  	 D_D 
R11          20  21      850
R5           22  3       100
QT14         24  18  2   Q_NPN 0.1
R21          6   2       2.67K
R20          3   6       13.08K
DZ2          25  26      D_5V1 
R19          1   26      16K
R18          14  3       250M
R17          25  14      380
R15          25  15      1.62K
QT16         1   20  15  Q_NPN 1
QT15         2   24  21  Q_PNP 0.1 
*OFF
R14          21  24      4K
C1           27  24      20P
R13          19  2       4K
QT13         24  27  18  Q_NPN 0.1
QT12         20  25  22  Q_NPN 1 
*OFF
QT11         20  28  2   Q_NPN 0.1
*OFF
QT10         20  11  1   Q_PNP 0.1
R10          17  27      16.5K
R9           5   4       1.9K
R8           4   23      26
R7           10  2       1.2K
R6           29  2       1K
QT9          11  11  1   Q_PNP 0.1
QT8          27  16  29  Q_NPN 0.1
QT4          15  6   17  Q_NPN 0.1
DZ1          2   9       D_5V6
R4           1   9       80K
R3           28  2       830
R2           13  28      4.97K
R1           8   13      7K

.MODEL D_5V1 D( IS=10F N=1.16 BV=5.1 IBV=0.5M CJO = 1P TT = 10p )
.MODEL D_5V6 D( IS=10F N=1.16 BV=5.6 IBV=5U CJO = 1P TT = 10p )
.MODEL Q_NPN NPN( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+       TF=10P TR=1N )
.MODEL Q_PNP PNP( IS=10F NF=1.16 NR=1.16 BF=80 CJC=1P CJE=2P  
+      TF=10P TR=1N )
.MODEL D_D D( IS=1F N=1.16 CJO = 1P TT = 10p )

.ENDS LM7824C




* Identical.

.SUBCKT LM7905-2  1    2    3            

DD4           4   5   D_6V3_0 
DD2           6   2   D_3V9_0 
DD1           7   2   D_4V7_0 
DD3           8   3   D_6V3_0 
C2            9  10  5P
C1            2   9  15P
QTU15         10   9   3   Q_PNP_0 1.000
R17          11  12  4.2K
QTU22          3  10  13   Q_NPN_0 3.000
R18           8   5  15.65K
R20          13  14  1K
R19           4  14  75
QTU31         12  11   4   Q_NPN_1 1.000
R16          15   1  160
R24          16   1  1.8K
C3           17   1  10P
QTU30         18  12  15   Q_NPN_1 1.000
QTU29         10  16   1   Q_NPN_1 1.000
R15          19   1  400
QTU28         10  20  19   Q_NPN_1 1.000
R14          21   1  200
QTU27         17  20  21   Q_NPN_1 1.000
R11          22  23  1K
R10          24  25  1K
QTU19         18  27  26   Q_NPN_1 1.000
R9            2  18  7.1K
QTU8          16  18   2   Q_PNP_0 1.000
QTU7          28  18   2   Q_PNP_0 1.000
QTU6          18  18   2   Q_PNP_0 1.000
QTU5          11  29   2   Q_PNP_0 1.000
QTU4          20  29   2   Q_PNP_0 1.000
QTU3           1  29   2   Q_PNP_0 1.000
QTU2           1  29   2   Q_PNP_0 1.000
R13          28   1  400
R12          30   1  400
QTU18         29  29  31   Q_NPN_1 1.000
QTU1          29  29   2   Q_PNP_0 1.000
R6           31  32  6.5K
R7           32  27  5.6K
R8           27  26  950
QTU10         33   6  26   Q_PNP_0 1.000
QTU17         34  35  33   Q_PNP_0 1.000
R5           36   1  2K
QTU24         34  34  36   Q_NPN_1 1.000
R1           37   6  6.3K
R2           37  38  670
R3           38  35  550
QTU9          38  35   6   Q_PNP_0 1.000
R4           39   1  2K
QTU23         35  34  39   Q_NPN_1 1.000
QTU16          1   7  35   Q_PNP_0 1.000
JT1           7   1   1  J_2N3458_N 
QTU14          3  17  23   Q_PNP_0 1.000
QTU13         17  17  23   Q_PNP_0 1.000
QTU12         17  17  25   Q_PNP_0 1.000
QTU11          9  17  25   Q_PNP_0 1.000
QTU32          3  13  14   Q_NPN_2 10.000
QTU26          9  20  28   Q_NPN_1 1.000
QTU25         20  20  30   Q_NPN_1 1.000
QTU21          2  40  22   Q_NPN_1 1.000
QTU20          2  37  24   Q_NPN_1 1.000
R21           2  40  4.29K
R22          40   3  500
R23          14   1  500M

.MODEL J_2N3458_N NJF( VTO=-3.05 BETA=699.53U LAMBDA=6M RD=1 RS=1 
+      CGD=2.81P CGS=2.91P M=227.1M PB=500M IS=114.41F 
+      VTOTC=-2.5M BETATCE=-500M KF=0 AF=1 )
.MODEL D_6V3_0  D( IS=10F N=1.24 BV=6.3 IBV=1M CJ0 = 1P TT = 10p )
.MODEL D_3V9_0  D( IS=10F N=1.24 BV=3.9 IBV=1M CJ0 = 1P TT = 10p )
.MODEL D_4V7_0  D( IS=10F N=1.24 BV=4.7 IBV=1M CJ0 = 1P TT = 10p )
.MODEL Q_PNP_0  PNP( IS=10F NF=1.04 NR=1.04 BF=50 CJC=1P CJE=2P
+      TF=10P TR=1N VAF=45)
.MODEL Q_NPN_0  NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.MODEL Q_NPN_1  NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.MODEL Q_NPN_2  NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.ENDS LM7905-2

* Identical but PIN 2 is now ADJUST instead of GND.
* LM117 seems to be the same model.

.SUBCKT LM317-1    1    2    3
D4            4   3  D_Z6V0
D3            5   6  D_Z6V3
D2            7   1  D_Z6V3
D1            3   8  D_Z6V3
QT26          1  10   9  Q_NPN 20.0
QT25          1  11  10  Q_NPN 2.0
QT24_2       13  12   5  Q_NPN 0.1
QT24         13  12  14  Q_NPN 0.1
QT23         17  16  15  Q_NPN 1.0
QT21         19  18   3  Q_NPN 0.1
QT19         21   3  20  Q_NPN 1.0
QT17         23   3  22  Q_NPN 0.1
QT13          1  25  24  Q_NPN 0.1
QT11         16  27  26  Q_NPN 0.1
QT7          30  29  28  Q_NPN 0.1
QT5          29  31   3  Q_NPN 0.1
QT3          33  31  32  Q_NPN 0.1
QT22_2       17  17   1  Q_PNP 1.0
QT22         16  17   1  Q_PNP 1.0
QT20          3  19  16  Q_PNP 0.1
QT18         21  21  16  Q_PNP 0.1
QT16         23  21  16  Q_PNP 0.1
QT15          3  23  25  Q_PNP 0.1
QT12          3  24  16  Q_PNP 0.1
QT9          27  30  34  Q_PNP 0.1
QT6           3  29  34  Q_PNP 0.1
QT14         25  33  35  Q_PNP 0.1
QT10         16  33  36  Q_PNP 0.1
QT8          34  33  37  Q_PNP 0.1
QT4          31  33  38  Q_PNP 0.1
QT2          33  33  39  Q_PNP 0.1
R27           4   2  50
R26           9   3  100M
R25           9  14  2
R24           5  14  160
R23           7   6  18K
R22          10   3  160
R21          12  13  400
R20          18  13  13K
R19          16  11  370
R18          15  10  130
R17          16  12  12K
C3           19  18  5P
R16          16  19  6.7K
R15          20  22  2.4K
R14          22   4  12K
C2           23   4  30P
C1           23   3  30P
R13          24   3  5.1K
R12          26   3  72
R11          27   3  5.8K
R10          28   3  4.1K
R9           32   3  180
R8           34  30  12.4K
R7           31  29  130
R6            8  31  100K
R5            1  35  5.6K
R4            1  36  82
R3            1  37  190
R2            1  38  310
R1            1  39  310
JT1           1   3   8  J_N

.MODEL D_Z6V0 D( IS=10F N=1.04 BV=6.0 IBV=1M CJ0 = 1P TT = 10p )
.MODEL D_Z6V3 D( IS=10F N=1.04 BV=6.3 IBV=1M CJ0 = 1P TT = 10p )
.MODEL Q_NPN NPN( IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P
+       TF=10P TR=1N VAF=90)
.MODEL Q_PNP PNP( IS=10F NF=1.04 NR=1.04 BF=50 CJC=1P CJE=2P
+      TF=10P TR=1N VAF=45)
.MODEL J_N NJF( VTO=-7 )

.ENDS LM317-1


.SUBCKT LM317-TI 1 2 3
J1 1 3 4 JN
Q2 5 5 6 QPL .1
Q3 5 8 9 QNL .2
Q4 8 5 7 QPL .1
Q5 81 8 3 QNL .2
Q6 3 81 10 QPL .2
Q7 12 81 13 QNL .2
Q8 10 5 11 QPL .2
Q9 14 12 10 QPL .2
Q10 16 5 17 QPL .2
Q11 16 14 15 QNL .2
Q12 3 20 16 QPL .2
Q13 1 19 20 QNL .2
Q14 19 5 18 QPL .2
Q15 3 21 19 QPL .2
Q16 21 22 16 QPL .2
Q17 21 3 24 QNL .2
Q18 22 22 16 QPL .2
Q19 22 3 241 QNL 2
Q20 3 25 16 QPL .2
Q21 25 26 3 QNL .2
Q22A 35 35 1 QPL 2
Q22B 16 35 1 QPL 2
Q23 35 16 30 QNL 2
Q24A 27 40 29 QNL .2
Q24B 27 40 28 QNL .2
Q25 1 31 41 QNL 5
Q26 1 41 32 QNL 50
D1 3 4 DZ
D2 33 1 DZ
D3 29 34 DZ
R1 1 6 310
R2 1 7 310
R3 1 11 190
R4 1 17 82
R5 1 18 5.6K
R6 4 8 100K
R7 8 81 130
R8 10 12 12.4K
R9 9 3 180
R10 13 3 4.1K
R11 14 3 5.8K
R12 15 3 72
R13 20 3 5.1K
R14 2 24 12K
R15 24 241 2.4K
R16 16 25 6.7K
R17 16 40 12K
R18 30 41 130
R19 16 31 370
R20 26 27 13K
R21 27 40 400
R22 3 41 160
R23 33 34 18K
R24 28 29 160
R25 28 32 3
R26 32 3 .1
C1 21 3 30PF
C2 21 2 30PF
C3 25 26 5PF
CBS1 5 3 2PF
CBS2 35 3 1PF
CBS3 22 3 1PF
.MODEL JN NJF(BETA=1E-4 VTO=-7)
.MODEL DZ D(BV=6.3)
.MODEL QNL NPN(EG=1.22 BF=80 RB=100 CCS=1.5PF TF=.3NS TR=6NS CJE=2PF
+ CJC=1PF VAF=100)
.MODEL QPL PNP(BF=40 RB=20 TF=.6NS TR=10NS CJE=1.5PF CJC=1PF VAF=50)
.ENDS LM317-TI



* LM317MOT Voltage Reg. (Motorola)

.SUBCKT LM317-MOT 1      2    3
*Connections  Input  Adj. Output
*LM317A voltage regulator - Motorola
J1 1 3 4 JN
Q2 5 5 6 QPL .1
Q3 5 8 9 QNL  .2
Q4 8 5 7 QPL .1
Q5 81 8 3 QNL .2
Q6 3 81 10 QPL .2
Q7 12 81 13 QNL  .2
Q8 10 5 11 QPL  .2 
Q9 14 12 10 QPL .2
Q10 16 5 17 QPL  .2
Q11 16 14 15 QNL .2
Q12 3 20 16 QPL .2
Q13 1 19 20 QNL .2
Q14 19 5 18 QPL .2
Q15 3 21 19 QPL .2
Q16 21 22 16 QPL .2
Q17 21 3 24 QNL   .2
Q18 22 22 16 QPL .2
Q19 22 3 241 QNL 2
Q20 3 25 16 QPL .2
Q21 25 26 3 QNL .2
Q22A 35 35 1 QPL 2
Q22B 16 35 1 QPL 2
Q23 35 16 30 QNL  2
Q24A 27 40 29 QNL .2
Q24B 27 40 28 QNL .2
Q25 1 31 41 QNL 5
Q26 1 41 32 QNL 50
D1 3 4 DZ
D2 33 1 DZ
D3 29 34 DZ
R1 1 6 310
R2 1 7 310
R3 1 11 230
R4 1 17 120
R5 1 18 5.6K
R6 4 8 125K
R7 8 81 135
R8 10 12 12.4K
R9 9 3 190
R10 13 3 3.6K
R11 14 3 5.8K
R12 15 3 110
R13 20 3 5.1K
R14 2 24 12.5K
R15 24 241 2.4K
R16 16 25 6.7K
R17 16 40 12K
R18 30 41 160
R19 16 31 170
R20 26 27 6.8K
R21 27 40 510
R22 3 41 200
R23 33 34 13K
R24 28 29 105
R25 28 32 4
R26 32 3 .1
C1 21 3 30PF
C2 21 2 30PF
C3 25 26 5PF
CBS1 5 3 2PF
CBS2 35 3 1PF
CBS3 22 3 1PF
.MODEL JN NJF(BETA=1E-4 VTO=-7)
.MODEL DZ D(BV=6.3)
.MODEL QNL NPN(EG=1.22 BF=80 RB=100 CCS=1.5PF TF=.3NS TR=6NS CJE=2PF
+ CJC=1PF VAF=100)
.MODEL QPL PNP(BF=40 RB=20 TF=.6NS TR=10NS CJE=1.5PF CJC=1PF VAF=50)
.ENDS LM317-MOT

*

*LM317 Voltage Reg. (Texas Inst)

.SUBCKT LM317-TI2 1      2    3
*Connections  Input  Adj. Output
*LM317 voltage regulator - Texas Instruments
J1 1 3 4 JN
Q2 5 5 6 QPL .1
Q3 5 8 9 QNL  .2
Q4 8 5 7 QPL .1
Q5 81 8 3 QNL .2
Q6 3 81 10 QPL .2
Q7 12 81 13 QNL  .2
Q8 10 5 11 QPL  .2 
Q9 14 12 10 QPL .2
Q10 16 5 17 QPL  .2
Q11 16 14 15 QNL .2
Q12 3 20 16 QPL .2
Q13 1 19 20 QNL .2
Q14 19 5 18 QPL .2
Q15 3 21 19 QPL .2
Q16 21 22 16 QPL .2
Q17 21 3 24 QNL   .2
Q18 22 22 16 QPL .2
Q19 22 3 241 QNL 2
Q20 3 25 16 QPL .2
Q21 25 26 3 QNL .2
Q22A 35 35 1 QPL 2
Q22B 16 35 1 QPL 2
Q23 35 16 30 QNL  2
Q24A 27 40 29 QNL .2
Q24B 27 40 28 QNL .2
Q25 1 31 41 QNL 5
Q26 1 41 32 QNL 50
D1 3 4 DZ
D2 33 1 DZ
D3 29 34 DZ
R1 1 6 310
R2 1 7 310
R3 1 11 190
R4 1 17 82
R5 1 18 5.6K
R6 4 8 100K
R7 8 81 130
R8 10 12 12.4K
R9 9 3 180
R10 13 3 4.1K
R11 14 3 5.8K
R12 15 3 72
R13 20 3 5.1K
R14 2 24 12K
R15 24 241 2.4K
R16 16 25 6.7K
R17 16 40 12K
R18 30 41 130
R19 16 31 370
R20 26 27 13K
R21 27 40 400
R22 3 41 160
R23 33 34 18K
R24 28 29 160
R25 28 32 3
R26 32 3 .1
C1 21 3 30PF
C2 21 2 30PF
C3 25 26 5PF
CBS1 5 3 2PF
CBS2 35 3 1PF
CBS3 22 3 1PF
.MODEL JN NJF(BETA=1E-4 VTO=-7)
.MODEL DZ D(BV=6.3)
.MODEL QNL NPN(EG=1.22 BF=80 RB=100 CCS=1.5PF TF=.3NS TR=6NS CJE=2PF
+ CJC=1PF VAF=100)
.MODEL QPL PNP(BF=40 RB=20 TF=.6NS TR=10NS CJE=1.5PF CJC=1PF VAF=50)
.ENDS LM317-TI2

*

*LM317 Voltage Reg. (Motorola)
.SUBCKT LM317-MOT2  1     2     3
*Connections     Input  Adj. Output
*LM317 voltage regulator
J1 1 3 4 JN 
Q2 5 5 6 QPL .25   
Q3 5 8 9 QNL    
Q4 8 5 7 QPL .25   
Q5 81 8 3 QNL   
Q6 3 81 10 QPL  
Q7 12 81 13 QNL 
Q8 10 5 11 QPL  
Q9 14 12 10 QPL 
Q10 16 5 17 QPL 
Q11 16 14 15 QNL
Q12 3 20 16 QPL 
Q13 1 19 20 QNL 
Q14 19 5 18 QPL 
Q15 3 21 19 QPL 
Q16 21 22 16 QPL
Q17 21 3 24 QNL 
Q18 22 22 16 QPL
Q19 22 3 241 QNL 10 
Q20 3 25 16 QPL 
Q21 25 26 3 QNL 
Q22A 35 35 1 QPL 2  
Q22B 16 35 1 QPL 2 
Q23 35 16 30 QNL 2 
Q24A 27 40 29 QNL   
Q24B 27 40 28 QNL   
Q25 1 31 41 QNL 40  
Q26 1 41 32 QNL 200 
D1 3 4 DZ   
D2 33 1 DZ  
D3 29 34 DZ 
R1 1 6 310  
R2 1 7 310  
R3 1 11 190 
R4 1 17 82  
R5 1 18 5.6K    
R6 4 8 125K 
R7 8 81 130 
R8 10 12 12.4K  
R9 9 3 180  
R10 13 3 4.1K   
R11 14 3 5.8K   
R12 15 3 72 
R13 20 3 5.1K   
R14 2 24 12K    
R15 24 241 2.4K 
R16 16 25 6.7K  
R17 16 40 12K   
R18 30 41 160   
R19 16 31 170   
R20 26 27 13K   
R21 27 40 400   
R22 3 41 160    
R23 33 34 18K   
R24 28 29 160   
R25 28 32 3 
R26 32 3 .1 
C1 21 3 30PF    
C2 21 2 30PF    
C3 25 26 5PF    
.MODEL JN NJF(BETA=1E-4 VTO=-7) 
.MODEL DZ D(BV=6.3) 
.MODEL QNL NPN(EG=1.22 BF=80 RB=100 CCS=2PF TF=.3NS TR=6NS CJE=3PF  
+ CJC=2PF VAF=100)   
.MODEL QPL PNP(BF=40 RB=20 TF=1NS TR=20NS CJE=6PF CJC=4PF VAF=100)   
.ENDS   LM317-MOT2


* from http://www.diyaudio.com/forums/showthread.php?threadid=5025
*LM337 negative voltage regulator
*Connections Input Adj. Output
.SUBCKT LM337-1 8 1 19
.MODEL QN NPN (BF=50 TF=1N CJC=1P)
.MODEL QPOUT PNP (BF=50 TF=1N RE=.2 CJC=1P)
.MODEL QP PNP CJC=1P TF=2N
.MODEL DN D
.MODEL D2 D BV=12 IBV=100U
R10 25 6 1K
Q3 8 17 16 QPOUT
Q4 8 25 17 QP
R18 19 17 250
R19 19 16 .3
G1 8 6 1 18 .1
C7 6 2 .04U
R24 2 8 100
I_ADJ 0 1 65U
R26 8 25 200K
Q5 25 4 19 QP
R27 16 4 200
R28 7 4 7K
D1 8 7 D2
D2 8 6 DN
V1 18 19 1.25
.ENDS


* modified from http://www.loutre.org/HIFI_LIB.LIB (quiescent current section biases to Input instead of Ground)
* MANUFACTURERS PART NO.= SG137A   (SILICON GENERAL)
* SUBTYPE: REGULATOR
* THIS FILE CONTAINS A PRE-RAD TEMPERATURE DEPENDENT MACROMODEL OF THE
* SG137A.
*
* PLEASE NOTE THE FOLLOWING:
*
* THIS MODEL CAN BE USED FROM -55 C TO 125 C WITH THE .TEMP
* STATEMENT.  IT INCLUDES POWER-UP AND POWER-DOWN EFFECTS.    IT IS
* NECESSARY TO SET ITL1=300  ITL2=300 WITH THE .OPTIONS COMMAND FOR 100%
* CONVERGENCE.  THESE  SETTINGS DETERMINE THE NUMBER OF ITERATIONS
* ALLOW FOR THE  CALCULATION OF THE DC AND BIAS PT VALUES WHEN THE
* STARTING POINT  IS CONSIDERED "BLIND" OR AN "EDUCATED GUESS".
* OTHER SETTINGS MAY WORK, BUT HAVE NOT BEEN TESTED YET.
*
* RIPPLE REJECTION, OUTPUT IMPEDANCE, QUIESCENT CURRENT, LINE
* TRANSIENT, DROPOUT, AND LOAD TRANSIENT RESPONSE ARE MODELED BASED
* ON LABORATORY MEASUREMENTS.  THE CORRELATION IS QUITE GOOD.
* CURRENT LIMITING AND ADJUSTMENT CURRENT BASED ON DATA SHEET
* INFORMATION ARE MODELED ACCURATELY.
*
*
*------------------------------------------------------------------
*
*
*
.SUBCKT LM337-2  3  1   2 
*                |  |   | 
*               IN  |   | 
*                  ADJ  |
*                      OUT  
*                       
*** VOLTAGE REFERENCE SECTION ***
LR 1 4  0.2709 TC1 = 7.8864E-4 TC2 = -2.8391E-5

RR 4 5 98.2994 TC=-0.0063, 6.2251E-5
CR 1 6 3P
RCR 6 7 150K
DZR 7 5 DZR
.MODEL DZR D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0.1P
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1.25
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 0.0001
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 2.2444E-6
+       TBV2 = 6.5556E-8
+       TRS1 = 0
+       TRS2 = 0
+ )
RZR 7 5 1MEG
DZ1 8 7 DZ1
.MODEL DZ1 D(
+         IS = 1E-14
+         RS = 1
+          N = 1
+         TT = 0
+        CJO = 1P
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 0.0001
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = -0.002847
+       TBV2 = 3.4722E-6
+       TRS1 = 0
+       TRS2 = 0
+ )
RQ 8 3 1.7546MEG TC=4.5212E-4,5.6515E-6
*** QUIESCENT CURRENT SECTION ***
FQ  1 3 VQ1 0.0625M
EQ1 24 3 1 7 1
VQ1 24 25 DC 0
RQ1 25 3 1 TC=-3.9528E-4,-1.1597E-5
*** ERROR AMPLIFIER ***
RIN 7 23 100K
E1  11 3 23 7 600
ROE1 9 11 10
D+ 9 13 DC
V+ 14 3 -1
E+ 13 14 1 3 1
.MODEL DC D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 10P
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
D- 12 9 DC
V- 12 3 DC 1
RP 9 10 151
CP 10 3 0.01U
E2 15 3 10 3 1
***
RB1 15 16 50
RB2 16 19 500 TC=-1.9327E-4,3.3434E-6
*** SHORT CIRCUIT AND FOLDBACK CURRENT SECTION ***
DSC 16 17 DMOD
ESC 17 3 POLY(1),(2,3) 2.447 -0.01
DFB 16 18 DMOD
EFB 18 3 POLY(1),(2,3) 12.5955 -1.2275 0.0457 -5.9169E-4
***
QP 20 19 3 QMOD
.MODEL QMOD NPN(
+         IS = 1E-14
+         BF = 500
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
*** DROPOUT VOLTAGE SECTION ***
RDO 23 22 0.1
DDO1 22 21 DDO
DDO2 21 20 DDO
.MODEL DDO D(
+         IS = 1E-14
+         RS = 0
+          N = 0.9687
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
***
RO 23 2 0.0017 TC=-0.07894, 0.001136
DDIS 3 23 DDIS
.MODEL DDIS D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 1PF
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.MODEL DMOD D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.ENDS LM337
