* A dual opamp ngspice model
* file name: TL072-dual.lib
.subckt TL072c 1 2 3 4 5 6 7 8
.include tl072.cir
XA 3 2 8 4 1 TL072
XB 5 6 8 4 7 TL072
.ends