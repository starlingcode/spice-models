.subckt SSI2130 1 2 3 4 5 7 8 9 10 11 12 13 14 15 16 17 18 20 21 22 23 24 26 27 28 29 31 32
R1 1 0 1Meg
R2 2 0 100k
R3 3 0 100k
R4 4 0 50k
R5 5 0 50k
R7 7 0 1m
R8 8 0 1.5k
R9 9 0 50k
R10 10 0 50k
R11 11 0 50k
R12 12 0 50k
R13 13 0 50k
R14 14 8 1m
R15 15 16 1m
R17 17 0 1Meg
R18 18 0 1Meg
R19 19 0 1Meg
R20 20 0 100k
R21 21 0 1m
R22 22 0 1m
R23 23 0 1Meg
R24 24 0 1Meg
R26 26 23 .1
R27 27 0 1.5k
R28 28 0 1Meg
R29 29 0 1Meg
R31 31 0 1Meg
R32 32 0 1Meg
.ends

