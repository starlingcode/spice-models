.subckt TRS_NORMAL 1 2 3
R1 1 2 .001
.ends

.subckt TRS_NORMAL_FAKE 1 2 3
R1 1 2 10Meg
.ends