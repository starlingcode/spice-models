**************** Discrete Diode Electrical Parameter ****************
* Product: MB2S
* Package: SOIC-4
* Bridge Rectifier 
* -------------------------------------------------------------------
.MODEL MB2SD D
+ n = 2.15337 is = 8.70529E-008 rs = 0.0464093 eg = 1.02043 xti = 3.0254
+ cjo = 2.36617E-011 vj = 0.866392 m = 0.324665 fc = 0.5 tt = 2.88539E-006 bv = 600
+ ibv = 0.0022 kf = 0 af = 1 t_measured = 27
* -------------------------------------------------------------------
* Creation: May-26-2009   Rev: 0.0
* Fairchild Semiconductor
.subckt MB2S 1 2 3 4
D1 1 3 MB2SD
D2 4 1 MB2SD
D3 4 2 MB2SD
D4 2 3 MB2SD
.ends