.subckt DG403 1 3 4 5 6 8 9 10 11 12 13 14 15 16
E1 i15 0 vol = '5.0 - V(15)'
S1 1 16 15 0 DGSWITCH
S2 3 4 i15 0 DGSWITCH
E2 i10 0 vol = '5.0 - V(10)'
S3 9 8 10 0 DGSWITCH
S4 5 6 i10 0 DGSWITCH
.model DGSWITCH SW (VT=3 VH=0 RON=30 ROFF=1e6)
.ends DG403