.include BLUE_LED.lib
.include RED_LED.lib
.subckt RB_BICOLOR 1 2
D1 1 2 BLUE_LED
D2 2 1 RED_LED
.ends