* A dual opamp ngspice model
* file name: TL072-dual.lib
.subckt TL074c 1 2 3 4 5 6 7 8 9 10 11 12 13 14
.include TL072.301
XA 3 2 4 11 1 TL072
XB 5 6 4 11 7 TL072
XC 10 9 4 11 8 TL072
XD 12 13 4 11 14 TL072
.ends