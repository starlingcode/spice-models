*SRC=MMBT3906;DI_MMBT3906;BJTs PNP; Si;  40.0V  0.200A  257MHz   Diodes Inc. Transistor
.MODEL DI_MMBT3906  PNP (IS=20.3f NF=1.00 BF=192 VAF=114
+ IKF=60.7m ISE=12.9p NE=2.00 BR=4.00 NR=1.00
+ VAR=20.0 IKR=0.150 RE=1.16 RB=4.63 RC=0.463
+ XTB=1.5 CJE=7.60p VJE=1.10 MJE=0.500 CJC=6.52p VJC=0.300
+ MJC=0.300 TF=589p TR=98.4n EG=1.12 )