.SUBCKT TL431 7 11 6
*             K A FDBK
.MODEL DCLAMP D (IS=13.5N RS=25M N=1.59 
+ CJO=45P VJ=.75 M=.302 TT=50.4N BV=34V IBV=1MA)
*V1 1 6 2.495 ; used for fixed reference, replaced with EB1 Limiter
EB1 1 6 Value = { IF ( V(7,6)> 2.495, 2.495, V(7,6) ) }
R1 6 2 15.6
C1 2 6 .5U
R2 2 3 100
C2 3 4 .08U
R3 4 6 10
G2 6 8 3 6 1.73
D1 5 8 DCLAMP
D2 7 8 DCLAMP
V4 5 6 2
G1 6 2 1 11 0.11
.ENDS