.SUBCKT THONKY S R T
R1 T R 0
.ENDS